module kareem
(
    input a, b, 
    output out
);
    and(out, a, b);
endmodule